.SUBCKT OPAMP1 3 2 1
RIN 1 2 10MEG
EGAIN 3 0   1 2  100K
.ENDS

